`timescale 1ns/1ps

// programmable bidirectional connection
module intercon_gate(
  input  shift_clk,
  input  shift_en,
  input  shift_i,
  output shift_o,

  inout  a,
  inout  b);

  // logic

endmodule
