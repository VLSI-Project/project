`timescale 1ns/1ps

// 3-input lookup table
module lut3(
  input  shift_clk,
  input  shift_en,
  input  shift_i,
  output shift_o,  

  input  a,
  input  b,
  input  c,
  output y);

  // logic to shift data in/out
  // logic to generate y

endmodule
