`timescale 1ns/1ps

// neg or pos edge D flip-flop or latch with async set/reset
module flop(
  input  shift_clk,
  input  shift_en,
  input  shift_i,
  output shift_o,

  input  flop_clk,
  input  set,
  input  rst,

  input  d,
  output q);

  // logic

endmodule
